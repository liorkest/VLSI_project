/*------------------------------------------------------------------------------
 * File          : divider_test.sv
 * Project       : RTL
 * Author        : eplkls
 * Creation date : Nov 23, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module divider_test #() ();

endmodule