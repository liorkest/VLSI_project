/*------------------------------------------------------------------------------
 * File          : noise_estimation.sv
 * Project       : RTL
 * Author        : eplkls
 * Creation date : Dec 12, 2024
 * Description   : This module receives 
 * 						1. block statistics (mean&variation) 
 * 						2. pixel-by-pixel of block
 * 					and calculates the pixel according to Weiner filter formula, 
 * 					for {TOTAL_SAMPLES} cycles, and goes to IDLE state again.
 *------------------------------------------------------------------------------*/

module wiener_calc #(
	parameter DATA_WIDTH = 8,        // Width of input data
	parameter TOTAL_SAMPLES = 64    // Total number of samples per block (MUST be power of 2)
)(
	input logic                   clk,
	input logic                   rst_n,
	input logic                   stats_ready,
	input logic [2*DATA_WIDTH-1:0] mean_of_block, // added 
	input logic [2*DATA_WIDTH-1:0] variance_of_block,
	input logic [2*DATA_WIDTH-1:0] noise_variance,
	input logic [DATA_WIDTH-1:0]  data_in,	      // the current pixel channel value 0-255
	input logic [31:0]            blocks_per_frame,
	// outputs
	output logic  [DATA_WIDTH-1:0] data_out,
	output logic [31:0]            data_count // starting from 1 to TOTAL_SAMPLES
);

// divider inst
logic [4*DATA_WIDTH-1 : 0] a;
logic [4*DATA_WIDTH-1 : 0] b;
logic [4*DATA_WIDTH-1 : 0] quotient; // result of 16.0 / 16.0 fixed point division = 16.16 format
logic [4*DATA_WIDTH-1 : 0] remainder;
logic divide_by_0;
DW_div divider (.*);

// divider inputs 
assign a = (variance_of_block >= noise_variance) ? 32'(variance_of_block - noise_variance) << 2*DATA_WIDTH : 32'(noise_variance - variance_of_block) << 2*DATA_WIDTH; // adjust to fixed point
assign b = (variance_of_block == 0) ? 32'b1 : 32'(variance_of_block);

logic [3*DATA_WIDTH-1:0]  data_out_unclipped;
logic quotient_sign;
logic data_mean_diff_sign;
logic [DATA_WIDTH-1:0] abs_data_mean_diff;
assign quotient_sign = (variance_of_block >= noise_variance) ? 1'b1 : 1'b0; // 1 - positive, 0 - negative
assign data_mean_diff_sign = (data_in >= mean_of_block) ? 1'b1 : 1'b0;
assign abs_data_mean_diff = (data_mean_diff_sign) ? data_in - mean_of_block[DATA_WIDTH-1:0] : mean_of_block[DATA_WIDTH-1:0] -data_in;

typedef enum logic [2:0] {
	IDLE = 0,
	CALCULATE = 1
 } state_t;

state_t state, next_state;

always_ff @(posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		state <= IDLE;
	end else begin
		state <= next_state;
	end
end

always_comb begin
	case (state) 
		IDLE: begin
			if (stats_ready) begin
				next_state = CALCULATE;
			end else begin
				next_state = IDLE;
			end
		end
		CALCULATE: begin
			if (data_count == TOTAL_SAMPLES + 2) begin  // +2 due to delay by 1 cycle of data_out
				next_state = IDLE;
			end else begin
				next_state = CALCULATE;
			end
		end
		default: begin
			next_state = IDLE;
		end
	endcase
end


// Data processing logic
always_ff @(posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		data_count<= 0;
		data_out <= 0;
		data_out_unclipped <= 0;
	end else begin
		// clipping 0-255 range
		if (data_out_unclipped < 0) data_out <= 0; 
		else if (data_out_unclipped > 255) data_out <= 255; 
		else data_out <= data_out_unclipped[DATA_WIDTH-1:0];
		
		if (state == IDLE && !next_state == CALCULATE) begin
			data_count <= 0;
		end else if (state == CALCULATE || next_state == CALCULATE) begin  // [12.12.24 LK] I wrote "next_state == calculate ",  otherwise we miss first sample!
			if (data_count == TOTAL_SAMPLES + 1) begin // +1 due to delay by 1 cycle of data_out
				data_count <= 0;
			end else begin
				data_count <= data_count + 1;
				if (quotient_sign == data_mean_diff_sign) begin
					data_out_unclipped <= mean_of_block + ((quotient * abs_data_mean_diff) >> 16);
				end else begin
					data_out_unclipped <= mean_of_block - ((quotient * abs_data_mean_diff) >> 16);
				end
			end
		end
	end
end

endmodule




