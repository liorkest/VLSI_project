/*------------------------------------------------------------------------------
 * File          : pixel_mean.sv
 * Project       : RTL
 * Author        : eplkls
 * Creation date : Dec 19, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module pixel_mean #() ();

endmodule